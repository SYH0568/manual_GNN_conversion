`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input reset,
    input clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 2'b0;
    localparam ST_DL_DETECTED = 2'b1;
    localparam ST_DL_REPORT = 2'b10;

    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        origin = 'b0;
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [560:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "myproject.Block_proc_U0";
                end
                1 : begin
                    proc_path = "myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0";
                end
                2 : begin
                    proc_path = "myproject.clone_vec_ap_uint_16_edge_index_config_1_U0";
                end
                3 : begin
                    proc_path = "myproject.clone_vec_ap_uint_16_edge_index_config_2_U0";
                end
                4 : begin
                    proc_path = "myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0";
                end
                5 : begin
                    proc_path = "myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0";
                end
                6 : begin
                    proc_path = "myproject.edge_aggregate_U0";
                end
                7 : begin
                    proc_path = "myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0";
                end
                8 : begin
                    proc_path = "myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [560:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [560:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [360:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    1: begin
                        if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    2: begin
                        if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    4: begin
                        if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_0_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_1_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_2_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_3_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_4_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_5_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_6_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_7_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_8_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_9_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_10_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_11_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_12_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_13_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_14_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_15_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_16_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_17_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_18_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_19_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_20_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_21_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_22_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_23_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_24_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_25_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_26_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_27_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_28_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_29_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_30_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_31_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_32_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_33_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_34_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_35_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_36_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_37_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_38_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_39_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_40_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_41_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_42_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_43_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_44_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_45_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_46_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy1_47_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    7: begin
                        if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_0_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_1_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_2_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_3_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_4_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_5_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_6_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_7_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_8_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_9_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_10_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_11_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_12_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_13_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_14_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_15_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_16_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_17_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_18_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_19_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_20_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_21_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_22_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_23_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_24_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_25_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_26_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_27_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_28_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_29_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_30_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_31_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_32_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_33_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_34_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_35_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_36_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_37_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_38_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_39_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_40_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_41_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_42_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_43_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_44_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_45_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_46_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_read) begin
                            chan_path = "myproject.node_attr_cpy2_47_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    2: begin
                        if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_14_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_16_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_18_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_20_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_22_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_24_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_26_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_28_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_30_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy2_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    1: begin
                        if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    2: begin
                        if (~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_0_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_1_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_2_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_3_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_4_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_5_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_6_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_7_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_8_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_9_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_10_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_11_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_12_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_13_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_14_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_15_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_16_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_17_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_18_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_19_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_20_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_21_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_22_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_23_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_24_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_25_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_26_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_27_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_28_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_29_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_30_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_write) begin
                            chan_path = "myproject.edge_index_cpy1_31_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy3_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    8: begin
                        if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_14_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_16_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_18_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_20_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_22_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_24_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_26_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_28_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_30_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_read) begin
                            chan_path = "myproject.edge_index_cpy4_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_0_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_1_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_2_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_3_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_4_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_5_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_6_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_7_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_8_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_9_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_10_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_11_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_12_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_13_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_14_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_15_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_16_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_17_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_18_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_19_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_20_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_21_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_22_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_23_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_24_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_25_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_26_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_27_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_28_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_29_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_30_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_31_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_32_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_33_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_34_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_35_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_36_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_37_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_38_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_39_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_40_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_41_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_42_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_43_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_44_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_45_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_46_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy1_47_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    2: begin
                        if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_14_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_16_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_18_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_20_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_22_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_24_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_26_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_28_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_30_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy2_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_myproject.layer7_out_0_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_0_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_1_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_1_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_2_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_2_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_3_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_3_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_4_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_4_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_5_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_5_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_6_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_6_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_7_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_7_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_8_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_8_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_9_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_9_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_10_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_10_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_11_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_11_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_12_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_12_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_13_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_13_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_14_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_14_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_15_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_15_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_16_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_16_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_17_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_17_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_18_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_18_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_19_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_19_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_20_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_20_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_21_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_21_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_22_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_22_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_23_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_23_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_24_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_24_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_25_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_25_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_26_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_26_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_27_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_27_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_28_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_28_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_29_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_29_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_30_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_30_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_31_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_31_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_32_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_32_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_33_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_33_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_34_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_34_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_35_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_35_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_36_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_36_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_37_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_37_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_38_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_38_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_39_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_39_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_40_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_40_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_41_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_41_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_42_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_42_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_43_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_43_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_44_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_44_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_45_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_45_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_46_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_46_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_47_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_47_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_48_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_48_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_49_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_49_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_50_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_50_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_51_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_51_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_52_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_52_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_53_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_53_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_54_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_54_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_55_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_55_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_56_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_56_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_57_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_57_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_58_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_58_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_59_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_59_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_60_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_60_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_61_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_61_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_62_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_62_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_63_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_63_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    0: begin
                        if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                            chan_path = "";
                            if (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]))) begin
                                $display("//      Deadlocked by sync logic between input processes");
                                $display("//      Please increase channel depth");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_myproject.layer7_out_0_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_0_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_1_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_1_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_2_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_2_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_3_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_3_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_4_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_4_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_5_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_5_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_6_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_6_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_7_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_7_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_8_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_8_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_9_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_9_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_10_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_10_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_11_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_11_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_12_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_12_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_13_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_13_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_14_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_14_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_15_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_15_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_16_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_16_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_17_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_17_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_18_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_18_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_19_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_19_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_20_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_20_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_21_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_21_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_22_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_22_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_23_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_23_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_24_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_24_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_25_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_25_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_26_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_26_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_27_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_27_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_28_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_28_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_29_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_29_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_30_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_30_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_31_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_31_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_32_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_32_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_33_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_33_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_34_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_34_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_35_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_35_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_36_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_36_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_37_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_37_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_38_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_38_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_39_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_39_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_40_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_40_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_41_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_41_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_42_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_42_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_43_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_43_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_44_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_44_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_45_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_45_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_46_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_46_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_47_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_47_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_48_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_48_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_49_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_49_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_50_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_50_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_51_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_51_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_52_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_52_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_53_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_53_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_54_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_54_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_55_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_55_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_56_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_56_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_57_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_57_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_58_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_58_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_59_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_59_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_60_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_60_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_61_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_61_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_62_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_62_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_63_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_63_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy1_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    8: begin
                        if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_read) begin
                            chan_path = "myproject.layer7_out_cpy2_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy1_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    3: begin
                        if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy3_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    7: begin
                        if (~AESL_inst_myproject.layer9_out_0_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_0_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_0_V_U";
                            if (~AESL_inst_myproject.layer9_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_1_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_1_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_1_V_U";
                            if (~AESL_inst_myproject.layer9_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_2_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_2_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_2_V_U";
                            if (~AESL_inst_myproject.layer9_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_3_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_3_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_3_V_U";
                            if (~AESL_inst_myproject.layer9_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_4_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_4_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_4_V_U";
                            if (~AESL_inst_myproject.layer9_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_5_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_5_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_5_V_U";
                            if (~AESL_inst_myproject.layer9_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_6_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_6_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_6_V_U";
                            if (~AESL_inst_myproject.layer9_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_7_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_7_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_7_V_U";
                            if (~AESL_inst_myproject.layer9_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_8_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_8_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_8_V_U";
                            if (~AESL_inst_myproject.layer9_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_9_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_9_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_9_V_U";
                            if (~AESL_inst_myproject.layer9_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_10_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_10_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_10_V_U";
                            if (~AESL_inst_myproject.layer9_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_11_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_11_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_11_V_U";
                            if (~AESL_inst_myproject.layer9_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_12_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_12_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_12_V_U";
                            if (~AESL_inst_myproject.layer9_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_13_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_13_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_13_V_U";
                            if (~AESL_inst_myproject.layer9_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_14_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_14_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_14_V_U";
                            if (~AESL_inst_myproject.layer9_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_15_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_15_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_15_V_U";
                            if (~AESL_inst_myproject.layer9_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_16_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_16_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_16_V_U";
                            if (~AESL_inst_myproject.layer9_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_17_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_17_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_17_V_U";
                            if (~AESL_inst_myproject.layer9_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_18_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_18_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_18_V_U";
                            if (~AESL_inst_myproject.layer9_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_19_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_19_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_19_V_U";
                            if (~AESL_inst_myproject.layer9_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_20_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_20_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_20_V_U";
                            if (~AESL_inst_myproject.layer9_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_21_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_21_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_21_V_U";
                            if (~AESL_inst_myproject.layer9_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_22_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_22_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_22_V_U";
                            if (~AESL_inst_myproject.layer9_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_23_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_23_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_23_V_U";
                            if (~AESL_inst_myproject.layer9_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_24_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_24_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_24_V_U";
                            if (~AESL_inst_myproject.layer9_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_25_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_25_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_25_V_U";
                            if (~AESL_inst_myproject.layer9_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_26_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_26_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_26_V_U";
                            if (~AESL_inst_myproject.layer9_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_27_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_27_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_27_V_U";
                            if (~AESL_inst_myproject.layer9_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_28_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_28_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_28_V_U";
                            if (~AESL_inst_myproject.layer9_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_29_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_29_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_29_V_U";
                            if (~AESL_inst_myproject.layer9_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_30_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_30_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_30_V_U";
                            if (~AESL_inst_myproject.layer9_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_31_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_31_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_31_V_U";
                            if (~AESL_inst_myproject.layer9_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_32_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_32_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_32_V_U";
                            if (~AESL_inst_myproject.layer9_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_33_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_33_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_33_V_U";
                            if (~AESL_inst_myproject.layer9_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_34_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_34_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_34_V_U";
                            if (~AESL_inst_myproject.layer9_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_35_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_35_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_35_V_U";
                            if (~AESL_inst_myproject.layer9_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_36_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_36_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_36_V_U";
                            if (~AESL_inst_myproject.layer9_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_37_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_37_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_37_V_U";
                            if (~AESL_inst_myproject.layer9_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_38_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_38_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_38_V_U";
                            if (~AESL_inst_myproject.layer9_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_39_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_39_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_39_V_U";
                            if (~AESL_inst_myproject.layer9_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_40_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_40_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_40_V_U";
                            if (~AESL_inst_myproject.layer9_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_41_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_41_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_41_V_U";
                            if (~AESL_inst_myproject.layer9_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_42_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_42_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_42_V_U";
                            if (~AESL_inst_myproject.layer9_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_43_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_43_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_43_V_U";
                            if (~AESL_inst_myproject.layer9_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_44_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_44_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_44_V_U";
                            if (~AESL_inst_myproject.layer9_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_45_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_45_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_45_V_U";
                            if (~AESL_inst_myproject.layer9_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_46_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_46_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_46_V_U";
                            if (~AESL_inst_myproject.layer9_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_47_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_47_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_47_V_U";
                            if (~AESL_inst_myproject.layer9_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_48_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_48_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_48_V_U";
                            if (~AESL_inst_myproject.layer9_out_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_49_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_49_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_49_V_U";
                            if (~AESL_inst_myproject.layer9_out_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_50_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_50_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_50_V_U";
                            if (~AESL_inst_myproject.layer9_out_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_51_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_51_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_51_V_U";
                            if (~AESL_inst_myproject.layer9_out_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_52_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_52_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_52_V_U";
                            if (~AESL_inst_myproject.layer9_out_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_53_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_53_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_53_V_U";
                            if (~AESL_inst_myproject.layer9_out_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_54_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_54_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_54_V_U";
                            if (~AESL_inst_myproject.layer9_out_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_55_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_55_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_55_V_U";
                            if (~AESL_inst_myproject.layer9_out_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_56_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_56_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_56_V_U";
                            if (~AESL_inst_myproject.layer9_out_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_57_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_57_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_57_V_U";
                            if (~AESL_inst_myproject.layer9_out_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_58_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_58_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_58_V_U";
                            if (~AESL_inst_myproject.layer9_out_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_59_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_59_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_59_V_U";
                            if (~AESL_inst_myproject.layer9_out_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_60_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_60_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_60_V_U";
                            if (~AESL_inst_myproject.layer9_out_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_61_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_61_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_61_V_U";
                            if (~AESL_inst_myproject.layer9_out_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_62_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_62_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_62_V_U";
                            if (~AESL_inst_myproject.layer9_out_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_63_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_63_V_U.t_read) begin
                            chan_path = "myproject.layer9_out_63_V_U";
                            if (~AESL_inst_myproject.layer9_out_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_0_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_1_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_2_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_3_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_4_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_5_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_6_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_7_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_8_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_9_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_10_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_11_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_12_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_13_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_14_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_15_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_16_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_17_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_18_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_19_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_20_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_21_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_22_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_23_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_24_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_25_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_26_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_27_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_28_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_29_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_30_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_31_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_32_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_33_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_34_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_35_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_36_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_37_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_38_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_39_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_40_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_41_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_42_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_43_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_44_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_45_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_46_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_write) begin
                            chan_path = "myproject.node_attr_cpy2_47_V_U";
                            if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_myproject.layer9_out_0_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_0_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_0_V_U";
                            if (~AESL_inst_myproject.layer9_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_1_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_1_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_1_V_U";
                            if (~AESL_inst_myproject.layer9_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_2_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_2_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_2_V_U";
                            if (~AESL_inst_myproject.layer9_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_3_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_3_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_3_V_U";
                            if (~AESL_inst_myproject.layer9_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_4_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_4_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_4_V_U";
                            if (~AESL_inst_myproject.layer9_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_5_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_5_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_5_V_U";
                            if (~AESL_inst_myproject.layer9_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_6_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_6_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_6_V_U";
                            if (~AESL_inst_myproject.layer9_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_7_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_7_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_7_V_U";
                            if (~AESL_inst_myproject.layer9_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_8_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_8_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_8_V_U";
                            if (~AESL_inst_myproject.layer9_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_9_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_9_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_9_V_U";
                            if (~AESL_inst_myproject.layer9_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_10_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_10_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_10_V_U";
                            if (~AESL_inst_myproject.layer9_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_11_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_11_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_11_V_U";
                            if (~AESL_inst_myproject.layer9_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_12_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_12_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_12_V_U";
                            if (~AESL_inst_myproject.layer9_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_13_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_13_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_13_V_U";
                            if (~AESL_inst_myproject.layer9_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_14_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_14_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_14_V_U";
                            if (~AESL_inst_myproject.layer9_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_15_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_15_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_15_V_U";
                            if (~AESL_inst_myproject.layer9_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_16_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_16_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_16_V_U";
                            if (~AESL_inst_myproject.layer9_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_17_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_17_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_17_V_U";
                            if (~AESL_inst_myproject.layer9_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_18_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_18_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_18_V_U";
                            if (~AESL_inst_myproject.layer9_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_19_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_19_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_19_V_U";
                            if (~AESL_inst_myproject.layer9_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_20_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_20_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_20_V_U";
                            if (~AESL_inst_myproject.layer9_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_21_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_21_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_21_V_U";
                            if (~AESL_inst_myproject.layer9_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_22_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_22_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_22_V_U";
                            if (~AESL_inst_myproject.layer9_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_23_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_23_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_23_V_U";
                            if (~AESL_inst_myproject.layer9_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_24_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_24_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_24_V_U";
                            if (~AESL_inst_myproject.layer9_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_25_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_25_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_25_V_U";
                            if (~AESL_inst_myproject.layer9_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_26_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_26_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_26_V_U";
                            if (~AESL_inst_myproject.layer9_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_27_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_27_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_27_V_U";
                            if (~AESL_inst_myproject.layer9_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_28_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_28_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_28_V_U";
                            if (~AESL_inst_myproject.layer9_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_29_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_29_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_29_V_U";
                            if (~AESL_inst_myproject.layer9_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_30_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_30_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_30_V_U";
                            if (~AESL_inst_myproject.layer9_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_31_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_31_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_31_V_U";
                            if (~AESL_inst_myproject.layer9_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_32_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_32_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_32_V_U";
                            if (~AESL_inst_myproject.layer9_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_33_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_33_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_33_V_U";
                            if (~AESL_inst_myproject.layer9_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_34_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_34_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_34_V_U";
                            if (~AESL_inst_myproject.layer9_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_35_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_35_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_35_V_U";
                            if (~AESL_inst_myproject.layer9_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_36_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_36_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_36_V_U";
                            if (~AESL_inst_myproject.layer9_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_37_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_37_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_37_V_U";
                            if (~AESL_inst_myproject.layer9_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_38_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_38_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_38_V_U";
                            if (~AESL_inst_myproject.layer9_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_39_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_39_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_39_V_U";
                            if (~AESL_inst_myproject.layer9_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_40_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_40_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_40_V_U";
                            if (~AESL_inst_myproject.layer9_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_41_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_41_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_41_V_U";
                            if (~AESL_inst_myproject.layer9_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_42_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_42_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_42_V_U";
                            if (~AESL_inst_myproject.layer9_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_43_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_43_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_43_V_U";
                            if (~AESL_inst_myproject.layer9_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_44_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_44_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_44_V_U";
                            if (~AESL_inst_myproject.layer9_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_45_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_45_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_45_V_U";
                            if (~AESL_inst_myproject.layer9_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_46_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_46_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_46_V_U";
                            if (~AESL_inst_myproject.layer9_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_47_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_47_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_47_V_U";
                            if (~AESL_inst_myproject.layer9_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_48_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_48_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_48_V_U";
                            if (~AESL_inst_myproject.layer9_out_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_49_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_49_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_49_V_U";
                            if (~AESL_inst_myproject.layer9_out_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_50_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_50_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_50_V_U";
                            if (~AESL_inst_myproject.layer9_out_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_51_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_51_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_51_V_U";
                            if (~AESL_inst_myproject.layer9_out_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_52_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_52_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_52_V_U";
                            if (~AESL_inst_myproject.layer9_out_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_53_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_53_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_53_V_U";
                            if (~AESL_inst_myproject.layer9_out_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_54_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_54_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_54_V_U";
                            if (~AESL_inst_myproject.layer9_out_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_55_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_55_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_55_V_U";
                            if (~AESL_inst_myproject.layer9_out_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_56_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_56_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_56_V_U";
                            if (~AESL_inst_myproject.layer9_out_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_57_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_57_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_57_V_U";
                            if (~AESL_inst_myproject.layer9_out_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_58_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_58_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_58_V_U";
                            if (~AESL_inst_myproject.layer9_out_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_59_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_59_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_59_V_U";
                            if (~AESL_inst_myproject.layer9_out_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_60_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_60_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_60_V_U";
                            if (~AESL_inst_myproject.layer9_out_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_61_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_61_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_61_V_U";
                            if (~AESL_inst_myproject.layer9_out_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_62_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_62_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_62_V_U";
                            if (~AESL_inst_myproject.layer9_out_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer9_out_63_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_63_V_U.i_write) begin
                            chan_path = "myproject.layer9_out_63_V_U";
                            if (~AESL_inst_myproject.layer9_out_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer9_out_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    8: begin
                        if (~AESL_inst_myproject.layer10_out_0_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_0_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_0_V_U";
                            if (~AESL_inst_myproject.layer10_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_1_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_1_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_1_V_U";
                            if (~AESL_inst_myproject.layer10_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_2_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_2_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_2_V_U";
                            if (~AESL_inst_myproject.layer10_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_3_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_3_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_3_V_U";
                            if (~AESL_inst_myproject.layer10_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_4_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_4_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_4_V_U";
                            if (~AESL_inst_myproject.layer10_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_5_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_5_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_5_V_U";
                            if (~AESL_inst_myproject.layer10_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_6_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_6_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_6_V_U";
                            if (~AESL_inst_myproject.layer10_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_7_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_7_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_7_V_U";
                            if (~AESL_inst_myproject.layer10_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_8_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_8_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_8_V_U";
                            if (~AESL_inst_myproject.layer10_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_9_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_9_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_9_V_U";
                            if (~AESL_inst_myproject.layer10_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_10_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_10_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_10_V_U";
                            if (~AESL_inst_myproject.layer10_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_11_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_11_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_11_V_U";
                            if (~AESL_inst_myproject.layer10_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_12_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_12_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_12_V_U";
                            if (~AESL_inst_myproject.layer10_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_13_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_13_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_13_V_U";
                            if (~AESL_inst_myproject.layer10_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_14_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_14_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_14_V_U";
                            if (~AESL_inst_myproject.layer10_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_15_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_15_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_15_V_U";
                            if (~AESL_inst_myproject.layer10_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_16_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_16_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_16_V_U";
                            if (~AESL_inst_myproject.layer10_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_17_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_17_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_17_V_U";
                            if (~AESL_inst_myproject.layer10_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_18_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_18_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_18_V_U";
                            if (~AESL_inst_myproject.layer10_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_19_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_19_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_19_V_U";
                            if (~AESL_inst_myproject.layer10_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_20_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_20_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_20_V_U";
                            if (~AESL_inst_myproject.layer10_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_21_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_21_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_21_V_U";
                            if (~AESL_inst_myproject.layer10_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_22_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_22_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_22_V_U";
                            if (~AESL_inst_myproject.layer10_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_23_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_23_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_23_V_U";
                            if (~AESL_inst_myproject.layer10_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_24_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_24_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_24_V_U";
                            if (~AESL_inst_myproject.layer10_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_25_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_25_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_25_V_U";
                            if (~AESL_inst_myproject.layer10_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_26_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_26_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_26_V_U";
                            if (~AESL_inst_myproject.layer10_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_27_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_27_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_27_V_U";
                            if (~AESL_inst_myproject.layer10_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_28_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_28_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_28_V_U";
                            if (~AESL_inst_myproject.layer10_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_29_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_29_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_29_V_U";
                            if (~AESL_inst_myproject.layer10_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_30_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_30_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_30_V_U";
                            if (~AESL_inst_myproject.layer10_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_31_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_31_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_31_V_U";
                            if (~AESL_inst_myproject.layer10_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_32_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_32_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_32_V_U";
                            if (~AESL_inst_myproject.layer10_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_33_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_33_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_33_V_U";
                            if (~AESL_inst_myproject.layer10_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_34_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_34_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_34_V_U";
                            if (~AESL_inst_myproject.layer10_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_35_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_35_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_35_V_U";
                            if (~AESL_inst_myproject.layer10_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_36_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_36_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_36_V_U";
                            if (~AESL_inst_myproject.layer10_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_37_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_37_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_37_V_U";
                            if (~AESL_inst_myproject.layer10_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_38_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_38_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_38_V_U";
                            if (~AESL_inst_myproject.layer10_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_39_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_39_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_39_V_U";
                            if (~AESL_inst_myproject.layer10_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_40_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_40_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_40_V_U";
                            if (~AESL_inst_myproject.layer10_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_41_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_41_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_41_V_U";
                            if (~AESL_inst_myproject.layer10_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_42_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_42_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_42_V_U";
                            if (~AESL_inst_myproject.layer10_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_43_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_43_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_43_V_U";
                            if (~AESL_inst_myproject.layer10_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_44_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_44_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_44_V_U";
                            if (~AESL_inst_myproject.layer10_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_45_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_45_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_45_V_U";
                            if (~AESL_inst_myproject.layer10_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_46_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_46_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_46_V_U";
                            if (~AESL_inst_myproject.layer10_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_47_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_47_V_U.t_read) begin
                            chan_path = "myproject.layer10_out_47_V_U";
                            if (~AESL_inst_myproject.layer10_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_myproject.layer10_out_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_0_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_0_V_U";
                            if (~AESL_inst_myproject.layer10_out_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_1_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_1_V_U";
                            if (~AESL_inst_myproject.layer10_out_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_2_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_2_V_U";
                            if (~AESL_inst_myproject.layer10_out_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_3_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_3_V_U";
                            if (~AESL_inst_myproject.layer10_out_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_4_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_4_V_U";
                            if (~AESL_inst_myproject.layer10_out_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_5_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_5_V_U";
                            if (~AESL_inst_myproject.layer10_out_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_6_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_6_V_U";
                            if (~AESL_inst_myproject.layer10_out_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_7_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_7_V_U";
                            if (~AESL_inst_myproject.layer10_out_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_8_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_8_V_U";
                            if (~AESL_inst_myproject.layer10_out_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_9_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_9_V_U";
                            if (~AESL_inst_myproject.layer10_out_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_10_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_10_V_U";
                            if (~AESL_inst_myproject.layer10_out_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_11_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_11_V_U";
                            if (~AESL_inst_myproject.layer10_out_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_12_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_12_V_U";
                            if (~AESL_inst_myproject.layer10_out_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_13_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_13_V_U";
                            if (~AESL_inst_myproject.layer10_out_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_14_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_14_V_U";
                            if (~AESL_inst_myproject.layer10_out_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_15_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_15_V_U";
                            if (~AESL_inst_myproject.layer10_out_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_16_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_16_V_U";
                            if (~AESL_inst_myproject.layer10_out_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_17_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_17_V_U";
                            if (~AESL_inst_myproject.layer10_out_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_18_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_18_V_U";
                            if (~AESL_inst_myproject.layer10_out_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_19_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_19_V_U";
                            if (~AESL_inst_myproject.layer10_out_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_20_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_20_V_U";
                            if (~AESL_inst_myproject.layer10_out_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_21_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_21_V_U";
                            if (~AESL_inst_myproject.layer10_out_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_22_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_22_V_U";
                            if (~AESL_inst_myproject.layer10_out_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_23_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_23_V_U";
                            if (~AESL_inst_myproject.layer10_out_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_24_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_24_V_U";
                            if (~AESL_inst_myproject.layer10_out_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_25_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_25_V_U";
                            if (~AESL_inst_myproject.layer10_out_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_26_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_26_V_U";
                            if (~AESL_inst_myproject.layer10_out_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_27_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_27_V_U";
                            if (~AESL_inst_myproject.layer10_out_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_28_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_28_V_U";
                            if (~AESL_inst_myproject.layer10_out_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_29_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_29_V_U";
                            if (~AESL_inst_myproject.layer10_out_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_30_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_30_V_U";
                            if (~AESL_inst_myproject.layer10_out_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_31_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_31_V_U";
                            if (~AESL_inst_myproject.layer10_out_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_32_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_32_V_U";
                            if (~AESL_inst_myproject.layer10_out_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_33_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_33_V_U";
                            if (~AESL_inst_myproject.layer10_out_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_34_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_34_V_U";
                            if (~AESL_inst_myproject.layer10_out_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_35_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_35_V_U";
                            if (~AESL_inst_myproject.layer10_out_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_36_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_36_V_U";
                            if (~AESL_inst_myproject.layer10_out_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_37_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_37_V_U";
                            if (~AESL_inst_myproject.layer10_out_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_38_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_38_V_U";
                            if (~AESL_inst_myproject.layer10_out_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_39_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_39_V_U";
                            if (~AESL_inst_myproject.layer10_out_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_40_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_40_V_U";
                            if (~AESL_inst_myproject.layer10_out_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_41_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_41_V_U";
                            if (~AESL_inst_myproject.layer10_out_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_42_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_42_V_U";
                            if (~AESL_inst_myproject.layer10_out_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_43_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_43_V_U";
                            if (~AESL_inst_myproject.layer10_out_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_44_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_44_V_U";
                            if (~AESL_inst_myproject.layer10_out_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_45_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_45_V_U";
                            if (~AESL_inst_myproject.layer10_out_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_46_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_46_V_U";
                            if (~AESL_inst_myproject.layer10_out_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer10_out_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_47_V_U.i_write) begin
                            chan_path = "myproject.layer10_out_47_V_U";
                            if (~AESL_inst_myproject.layer10_out_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer10_out_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_0_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_1_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_2_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_3_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_4_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_5_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_6_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_7_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_8_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_9_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_10_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_11_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_12_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_13_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_14_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_15_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_16_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_17_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_18_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_19_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_20_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_21_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_22_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_23_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_24_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_25_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_26_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_27_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_28_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_29_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_30_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_31_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_32_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_33_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_34_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_35_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_36_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_37_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_38_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_39_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_40_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_41_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_42_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_43_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_44_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_45_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_46_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_47_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_48_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_49_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_50_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_51_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_52_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_53_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_54_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_55_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_56_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_57_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_58_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_59_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_60_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_61_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_62_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_write) begin
                            chan_path = "myproject.layer7_out_cpy2_63_V_U";
                            if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    3: begin
                        if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_0_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_1_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_2_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_3_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_4_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_5_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_6_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_7_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_8_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_9_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_10_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_11_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_12_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_13_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_14_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_15_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_16_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_17_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_18_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_19_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_20_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_21_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_22_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_23_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_24_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_25_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_26_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_27_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_28_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_29_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_30_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_write) begin
                            chan_path = "myproject.edge_index_cpy4_31_V_U";
                            if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        wait (reset == 1);
        cycle_id = 1;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end(cycle_id - 1);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
