`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [2:0] proc_dep_vld_vec_0;
    reg [2:0] proc_dep_vld_vec_0_reg;
    wire [2:0] in_chan_dep_vld_vec_0;
    wire [26:0] in_chan_dep_data_vec_0;
    wire [2:0] token_in_vec_0;
    wire [2:0] out_chan_dep_vld_vec_0;
    wire [8:0] out_chan_dep_data_0;
    wire [2:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [8:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [8:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_4_0;
    wire [8:0] dep_chan_data_4_0;
    wire token_4_0;
    wire [3:0] proc_dep_vld_vec_1;
    reg [3:0] proc_dep_vld_vec_1_reg;
    wire [3:0] in_chan_dep_vld_vec_1;
    wire [35:0] in_chan_dep_data_vec_1;
    wire [3:0] token_in_vec_1;
    wire [3:0] out_chan_dep_vld_vec_1;
    wire [8:0] out_chan_dep_data_1;
    wire [3:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [8:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [8:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_4_1;
    wire [8:0] dep_chan_data_4_1;
    wire token_4_1;
    wire dep_chan_vld_7_1;
    wire [8:0] dep_chan_data_7_1;
    wire token_7_1;
    wire [2:0] proc_dep_vld_vec_2;
    reg [2:0] proc_dep_vld_vec_2_reg;
    wire [3:0] in_chan_dep_vld_vec_2;
    wire [35:0] in_chan_dep_data_vec_2;
    wire [3:0] token_in_vec_2;
    wire [2:0] out_chan_dep_vld_vec_2;
    wire [8:0] out_chan_dep_data_2;
    wire [2:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [8:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [8:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [8:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_4_2;
    wire [8:0] dep_chan_data_4_2;
    wire token_4_2;
    wire [2:0] proc_dep_vld_vec_3;
    reg [2:0] proc_dep_vld_vec_3_reg;
    wire [1:0] in_chan_dep_vld_vec_3;
    wire [17:0] in_chan_dep_data_vec_3;
    wire [1:0] token_in_vec_3;
    wire [2:0] out_chan_dep_vld_vec_3;
    wire [8:0] out_chan_dep_data_3;
    wire [2:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_6_3;
    wire [8:0] dep_chan_data_6_3;
    wire token_6_3;
    wire dep_chan_vld_8_3;
    wire [8:0] dep_chan_data_8_3;
    wire token_8_3;
    wire [3:0] proc_dep_vld_vec_4;
    reg [3:0] proc_dep_vld_vec_4_reg;
    wire [3:0] in_chan_dep_vld_vec_4;
    wire [35:0] in_chan_dep_data_vec_4;
    wire [3:0] token_in_vec_4;
    wire [3:0] out_chan_dep_vld_vec_4;
    wire [8:0] out_chan_dep_data_4;
    wire [3:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_0_4;
    wire [8:0] dep_chan_data_0_4;
    wire token_0_4;
    wire dep_chan_vld_1_4;
    wire [8:0] dep_chan_data_1_4;
    wire token_1_4;
    wire dep_chan_vld_2_4;
    wire [8:0] dep_chan_data_2_4;
    wire token_2_4;
    wire dep_chan_vld_5_4;
    wire [8:0] dep_chan_data_5_4;
    wire token_5_4;
    wire [2:0] proc_dep_vld_vec_5;
    reg [2:0] proc_dep_vld_vec_5_reg;
    wire [2:0] in_chan_dep_vld_vec_5;
    wire [26:0] in_chan_dep_data_vec_5;
    wire [2:0] token_in_vec_5;
    wire [2:0] out_chan_dep_vld_vec_5;
    wire [8:0] out_chan_dep_data_5;
    wire [2:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_4_5;
    wire [8:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [8:0] dep_chan_data_6_5;
    wire token_6_5;
    wire dep_chan_vld_8_5;
    wire [8:0] dep_chan_data_8_5;
    wire token_8_5;
    wire [2:0] proc_dep_vld_vec_6;
    reg [2:0] proc_dep_vld_vec_6_reg;
    wire [2:0] in_chan_dep_vld_vec_6;
    wire [26:0] in_chan_dep_data_vec_6;
    wire [2:0] token_in_vec_6;
    wire [2:0] out_chan_dep_vld_vec_6;
    wire [8:0] out_chan_dep_data_6;
    wire [2:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_3_6;
    wire [8:0] dep_chan_data_3_6;
    wire token_3_6;
    wire dep_chan_vld_5_6;
    wire [8:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_7_6;
    wire [8:0] dep_chan_data_7_6;
    wire token_7_6;
    wire [2:0] proc_dep_vld_vec_7;
    reg [2:0] proc_dep_vld_vec_7_reg;
    wire [2:0] in_chan_dep_vld_vec_7;
    wire [26:0] in_chan_dep_data_vec_7;
    wire [2:0] token_in_vec_7;
    wire [2:0] out_chan_dep_vld_vec_7;
    wire [8:0] out_chan_dep_data_7;
    wire [2:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_1_7;
    wire [8:0] dep_chan_data_1_7;
    wire token_1_7;
    wire dep_chan_vld_6_7;
    wire [8:0] dep_chan_data_6_7;
    wire token_6_7;
    wire dep_chan_vld_8_7;
    wire [8:0] dep_chan_data_8_7;
    wire token_8_7;
    wire [2:0] proc_dep_vld_vec_8;
    reg [2:0] proc_dep_vld_vec_8_reg;
    wire [2:0] in_chan_dep_vld_vec_8;
    wire [26:0] in_chan_dep_data_vec_8;
    wire [2:0] token_in_vec_8;
    wire [2:0] out_chan_dep_vld_vec_8;
    wire [8:0] out_chan_dep_data_8;
    wire [2:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_3_8;
    wire [8:0] dep_chan_data_3_8;
    wire token_3_8;
    wire dep_chan_vld_5_8;
    wire [8:0] dep_chan_data_5_8;
    wire token_5_8;
    wire dep_chan_vld_7_8;
    wire [8:0] dep_chan_data_7_8;
    wire token_7_8;
    wire [8:0] dl_in_vec;
    wire dl_detect_out;
    wire [8:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done;
        end
    end

    reg ap_done_reg_2;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done;
        end
    end

    reg ap_done_reg_3;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done;
        end
    end

    reg ap_done_reg_4;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_4 <= 'b0;
        end
        else begin
            ap_done_reg_4 <= AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done;
        end
    end

    reg ap_done_reg_5;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_5 <= 'b0;
        end
        else begin
            ap_done_reg_5 <= AESL_inst_myproject.edge_aggregate_U0.ap_done;
        end
    end

    reg ap_done_reg_6;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_6 <= 'b0;
        end
        else begin
            ap_done_reg_6 <= AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done;
        end
    end

    reg ap_done_reg_7;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_7 <= 'b0;
        end
        else begin
            ap_done_reg_7 <= AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$Block_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$Block_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$Block_proc_U0$ap_idle <= AESL_inst_myproject.Block_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.Block_proc_U0
    AESL_deadlock_detect_unit #(9, 0, 3, 3) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (((AESL_inst_myproject.Block_proc_U0_ap_ready_count[0]) & AESL_inst_myproject.Block_proc_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[8 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[17 : 9] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_4_0;
    assign in_chan_dep_data_vec_0[26 : 18] = dep_chan_data_4_0;
    assign token_in_vec_0[2] = token_4_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[1];
    assign dep_chan_vld_0_4 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_4 = out_chan_dep_data_0;
    assign token_0_4 = token_out_vec_0[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0$ap_idle <= AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0
    AESL_deadlock_detect_unit #(9, 1, 4, 4) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_read | ((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_read | ~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_read);
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (((AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[8 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[17 : 9] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_4_1;
    assign in_chan_dep_data_vec_1[26 : 18] = dep_chan_data_4_1;
    assign token_in_vec_1[2] = token_4_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_7_1;
    assign in_chan_dep_data_vec_1[35 : 27] = dep_chan_data_7_1;
    assign token_in_vec_1[3] = token_7_1;
    assign dep_chan_vld_1_4 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_4 = out_chan_dep_data_1;
    assign token_1_4 = token_out_vec_1[0];
    assign dep_chan_vld_1_7 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_7 = out_chan_dep_data_1;
    assign token_1_7 = token_out_vec_1[1];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[2];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_1_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_1_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_1_U0$ap_idle <= AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0
    AESL_deadlock_detect_unit #(9, 2, 4, 3) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_read | ((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (((AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0]) & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[8 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[17 : 9] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[26 : 18] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_4_2;
    assign in_chan_dep_data_vec_2[35 : 27] = dep_chan_data_4_2;
    assign token_in_vec_2[3] = token_4_2;
    assign dep_chan_vld_2_4 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_4 = out_chan_dep_data_2;
    assign token_2_4 = token_out_vec_2[0];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[1];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_2_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_2_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$clone_vec_ap_uint_16_edge_index_config_2_U0$ap_idle <= AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0
    AESL_deadlock_detect_unit #(9, 3, 2, 3) AESL_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_0_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_1_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_2_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_3_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_4_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_5_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_6_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_7_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_8_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_9_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_10_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_11_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_12_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_13_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_14_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_15_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_16_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_17_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_18_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_19_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_20_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_21_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_22_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_23_12_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_24_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_25_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_26_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_27_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_28_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_29_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_30_11_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_0_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_1_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_2_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_3_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_4_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_5_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_6_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_7_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_8_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_9_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_10_V_U.if_write | ~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_empty_n & (AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy1_31_11_V_U.if_write);
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_read);
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_read | ~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_2_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_6_3;
    assign in_chan_dep_data_vec_3[8 : 0] = dep_chan_data_6_3;
    assign token_in_vec_3[0] = token_6_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_8_3;
    assign in_chan_dep_data_vec_3[17 : 9] = dep_chan_data_8_3;
    assign token_in_vec_3[1] = token_8_3;
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[0];
    assign dep_chan_vld_3_6 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_6 = out_chan_dep_data_3;
    assign token_3_6 = token_out_vec_3[1];
    assign dep_chan_vld_3_8 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_8 = out_chan_dep_data_3;
    assign token_3_8 = token_out_vec_3[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0$ap_idle <= AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0
    AESL_deadlock_detect_unit #(9, 4, 4, 4) AESL_deadlock_detect_unit_4 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (~AESL_inst_myproject.node_attr_cpy1_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_0_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_1_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_2_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_3_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_4_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_5_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_6_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_7_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_8_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_9_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_10_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_11_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_12_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_13_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_14_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_15_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_16_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_17_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_18_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_19_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_20_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_21_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_22_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_23_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_24_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_25_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_26_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_27_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_28_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_29_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_30_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_31_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_32_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_33_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_34_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_35_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_36_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_37_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_38_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_39_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_40_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_41_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_42_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_43_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_44_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_45_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_46_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy1_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy1_47_V_U.i_write | ((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_node_attr_config_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (~AESL_inst_myproject.edge_index_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_0_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_1_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_2_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_3_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_4_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_5_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_6_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_7_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_8_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_9_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_10_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_11_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_12_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_13_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_14_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_15_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_16_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_17_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_18_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_19_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_20_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_21_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_22_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_23_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_24_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_25_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_26_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_27_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_28_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_29_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_30_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy2_31_V_U.i_write | ((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.clone_vec_ap_uint_16_edge_index_config_1_U0_ap_ready_count[0])));
    assign proc_dep_vld_vec_4[2] = dl_detect_out ? proc_dep_vld_vec_4_reg[2] : (~AESL_inst_myproject.layer7_out_0_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_0_V_U.t_read | ~AESL_inst_myproject.layer7_out_1_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_1_V_U.t_read | ~AESL_inst_myproject.layer7_out_2_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_2_V_U.t_read | ~AESL_inst_myproject.layer7_out_3_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_3_V_U.t_read | ~AESL_inst_myproject.layer7_out_4_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_4_V_U.t_read | ~AESL_inst_myproject.layer7_out_5_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_5_V_U.t_read | ~AESL_inst_myproject.layer7_out_6_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_6_V_U.t_read | ~AESL_inst_myproject.layer7_out_7_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_7_V_U.t_read | ~AESL_inst_myproject.layer7_out_8_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_8_V_U.t_read | ~AESL_inst_myproject.layer7_out_9_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_9_V_U.t_read | ~AESL_inst_myproject.layer7_out_10_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_10_V_U.t_read | ~AESL_inst_myproject.layer7_out_11_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_11_V_U.t_read | ~AESL_inst_myproject.layer7_out_12_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_12_V_U.t_read | ~AESL_inst_myproject.layer7_out_13_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_13_V_U.t_read | ~AESL_inst_myproject.layer7_out_14_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_14_V_U.t_read | ~AESL_inst_myproject.layer7_out_15_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_15_V_U.t_read | ~AESL_inst_myproject.layer7_out_16_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_16_V_U.t_read | ~AESL_inst_myproject.layer7_out_17_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_17_V_U.t_read | ~AESL_inst_myproject.layer7_out_18_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_18_V_U.t_read | ~AESL_inst_myproject.layer7_out_19_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_19_V_U.t_read | ~AESL_inst_myproject.layer7_out_20_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_20_V_U.t_read | ~AESL_inst_myproject.layer7_out_21_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_21_V_U.t_read | ~AESL_inst_myproject.layer7_out_22_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_22_V_U.t_read | ~AESL_inst_myproject.layer7_out_23_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_23_V_U.t_read | ~AESL_inst_myproject.layer7_out_24_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_24_V_U.t_read | ~AESL_inst_myproject.layer7_out_25_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_25_V_U.t_read | ~AESL_inst_myproject.layer7_out_26_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_26_V_U.t_read | ~AESL_inst_myproject.layer7_out_27_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_27_V_U.t_read | ~AESL_inst_myproject.layer7_out_28_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_28_V_U.t_read | ~AESL_inst_myproject.layer7_out_29_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_29_V_U.t_read | ~AESL_inst_myproject.layer7_out_30_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_30_V_U.t_read | ~AESL_inst_myproject.layer7_out_31_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_31_V_U.t_read | ~AESL_inst_myproject.layer7_out_32_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_32_V_U.t_read | ~AESL_inst_myproject.layer7_out_33_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_33_V_U.t_read | ~AESL_inst_myproject.layer7_out_34_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_34_V_U.t_read | ~AESL_inst_myproject.layer7_out_35_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_35_V_U.t_read | ~AESL_inst_myproject.layer7_out_36_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_36_V_U.t_read | ~AESL_inst_myproject.layer7_out_37_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_37_V_U.t_read | ~AESL_inst_myproject.layer7_out_38_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_38_V_U.t_read | ~AESL_inst_myproject.layer7_out_39_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_39_V_U.t_read | ~AESL_inst_myproject.layer7_out_40_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_40_V_U.t_read | ~AESL_inst_myproject.layer7_out_41_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_41_V_U.t_read | ~AESL_inst_myproject.layer7_out_42_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_42_V_U.t_read | ~AESL_inst_myproject.layer7_out_43_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_43_V_U.t_read | ~AESL_inst_myproject.layer7_out_44_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_44_V_U.t_read | ~AESL_inst_myproject.layer7_out_45_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_45_V_U.t_read | ~AESL_inst_myproject.layer7_out_46_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_46_V_U.t_read | ~AESL_inst_myproject.layer7_out_47_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_47_V_U.t_read | ~AESL_inst_myproject.layer7_out_48_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_48_V_U.t_read | ~AESL_inst_myproject.layer7_out_49_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_49_V_U.t_read | ~AESL_inst_myproject.layer7_out_50_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_50_V_U.t_read | ~AESL_inst_myproject.layer7_out_51_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_51_V_U.t_read | ~AESL_inst_myproject.layer7_out_52_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_52_V_U.t_read | ~AESL_inst_myproject.layer7_out_53_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_53_V_U.t_read | ~AESL_inst_myproject.layer7_out_54_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_54_V_U.t_read | ~AESL_inst_myproject.layer7_out_55_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_55_V_U.t_read | ~AESL_inst_myproject.layer7_out_56_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_56_V_U.t_read | ~AESL_inst_myproject.layer7_out_57_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_57_V_U.t_read | ~AESL_inst_myproject.layer7_out_58_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_58_V_U.t_read | ~AESL_inst_myproject.layer7_out_59_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_59_V_U.t_read | ~AESL_inst_myproject.layer7_out_60_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_60_V_U.t_read | ~AESL_inst_myproject.layer7_out_61_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_61_V_U.t_read | ~AESL_inst_myproject.layer7_out_62_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_62_V_U.t_read | ~AESL_inst_myproject.layer7_out_63_V_U.i_full_n & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_done & deadlock_detector.ap_done_reg_3 & ~AESL_inst_myproject.layer7_out_63_V_U.t_read);
    assign proc_dep_vld_vec_4[3] = dl_detect_out ? proc_dep_vld_vec_4_reg[3] : (((AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0_ap_ready_count[0]) & AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config7_U0.ap_idle & ~(AESL_inst_myproject.Block_proc_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_0_4;
    assign in_chan_dep_data_vec_4[8 : 0] = dep_chan_data_0_4;
    assign token_in_vec_4[0] = token_0_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_1_4;
    assign in_chan_dep_data_vec_4[17 : 9] = dep_chan_data_1_4;
    assign token_in_vec_4[1] = token_1_4;
    assign in_chan_dep_vld_vec_4[2] = dep_chan_vld_2_4;
    assign in_chan_dep_data_vec_4[26 : 18] = dep_chan_data_2_4;
    assign token_in_vec_4[2] = token_2_4;
    assign in_chan_dep_vld_vec_4[3] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[35 : 27] = dep_chan_data_5_4;
    assign token_in_vec_4[3] = token_5_4;
    assign dep_chan_vld_4_1 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_1 = out_chan_dep_data_4;
    assign token_4_1 = token_out_vec_4[0];
    assign dep_chan_vld_4_2 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_2 = out_chan_dep_data_4;
    assign token_4_2 = token_out_vec_4[1];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[2];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[2];
    assign dep_chan_vld_4_0 = out_chan_dep_vld_vec_4[3];
    assign dep_chan_data_4_0 = out_chan_dep_data_4;
    assign token_4_0 = token_out_vec_4[3];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0$ap_idle <= AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0
    AESL_deadlock_detect_unit #(9, 5, 3, 3) AESL_deadlock_detect_unit_5 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (~AESL_inst_myproject.layer7_out_0_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_0_V_U.i_write | ~AESL_inst_myproject.layer7_out_1_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_1_V_U.i_write | ~AESL_inst_myproject.layer7_out_2_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_2_V_U.i_write | ~AESL_inst_myproject.layer7_out_3_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_3_V_U.i_write | ~AESL_inst_myproject.layer7_out_4_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_4_V_U.i_write | ~AESL_inst_myproject.layer7_out_5_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_5_V_U.i_write | ~AESL_inst_myproject.layer7_out_6_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_6_V_U.i_write | ~AESL_inst_myproject.layer7_out_7_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_7_V_U.i_write | ~AESL_inst_myproject.layer7_out_8_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_8_V_U.i_write | ~AESL_inst_myproject.layer7_out_9_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_9_V_U.i_write | ~AESL_inst_myproject.layer7_out_10_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_10_V_U.i_write | ~AESL_inst_myproject.layer7_out_11_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_11_V_U.i_write | ~AESL_inst_myproject.layer7_out_12_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_12_V_U.i_write | ~AESL_inst_myproject.layer7_out_13_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_13_V_U.i_write | ~AESL_inst_myproject.layer7_out_14_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_14_V_U.i_write | ~AESL_inst_myproject.layer7_out_15_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_15_V_U.i_write | ~AESL_inst_myproject.layer7_out_16_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_16_V_U.i_write | ~AESL_inst_myproject.layer7_out_17_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_17_V_U.i_write | ~AESL_inst_myproject.layer7_out_18_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_18_V_U.i_write | ~AESL_inst_myproject.layer7_out_19_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_19_V_U.i_write | ~AESL_inst_myproject.layer7_out_20_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_20_V_U.i_write | ~AESL_inst_myproject.layer7_out_21_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_21_V_U.i_write | ~AESL_inst_myproject.layer7_out_22_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_22_V_U.i_write | ~AESL_inst_myproject.layer7_out_23_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_23_V_U.i_write | ~AESL_inst_myproject.layer7_out_24_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_24_V_U.i_write | ~AESL_inst_myproject.layer7_out_25_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_25_V_U.i_write | ~AESL_inst_myproject.layer7_out_26_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_26_V_U.i_write | ~AESL_inst_myproject.layer7_out_27_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_27_V_U.i_write | ~AESL_inst_myproject.layer7_out_28_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_28_V_U.i_write | ~AESL_inst_myproject.layer7_out_29_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_29_V_U.i_write | ~AESL_inst_myproject.layer7_out_30_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_30_V_U.i_write | ~AESL_inst_myproject.layer7_out_31_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_31_V_U.i_write | ~AESL_inst_myproject.layer7_out_32_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_32_V_U.i_write | ~AESL_inst_myproject.layer7_out_33_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_33_V_U.i_write | ~AESL_inst_myproject.layer7_out_34_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_34_V_U.i_write | ~AESL_inst_myproject.layer7_out_35_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_35_V_U.i_write | ~AESL_inst_myproject.layer7_out_36_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_36_V_U.i_write | ~AESL_inst_myproject.layer7_out_37_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_37_V_U.i_write | ~AESL_inst_myproject.layer7_out_38_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_38_V_U.i_write | ~AESL_inst_myproject.layer7_out_39_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_39_V_U.i_write | ~AESL_inst_myproject.layer7_out_40_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_40_V_U.i_write | ~AESL_inst_myproject.layer7_out_41_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_41_V_U.i_write | ~AESL_inst_myproject.layer7_out_42_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_42_V_U.i_write | ~AESL_inst_myproject.layer7_out_43_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_43_V_U.i_write | ~AESL_inst_myproject.layer7_out_44_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_44_V_U.i_write | ~AESL_inst_myproject.layer7_out_45_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_45_V_U.i_write | ~AESL_inst_myproject.layer7_out_46_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_46_V_U.i_write | ~AESL_inst_myproject.layer7_out_47_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_47_V_U.i_write | ~AESL_inst_myproject.layer7_out_48_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_48_V_U.i_write | ~AESL_inst_myproject.layer7_out_49_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_49_V_U.i_write | ~AESL_inst_myproject.layer7_out_50_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_50_V_U.i_write | ~AESL_inst_myproject.layer7_out_51_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_51_V_U.i_write | ~AESL_inst_myproject.layer7_out_52_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_52_V_U.i_write | ~AESL_inst_myproject.layer7_out_53_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_53_V_U.i_write | ~AESL_inst_myproject.layer7_out_54_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_54_V_U.i_write | ~AESL_inst_myproject.layer7_out_55_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_55_V_U.i_write | ~AESL_inst_myproject.layer7_out_56_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_56_V_U.i_write | ~AESL_inst_myproject.layer7_out_57_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_57_V_U.i_write | ~AESL_inst_myproject.layer7_out_58_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_58_V_U.i_write | ~AESL_inst_myproject.layer7_out_59_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_59_V_U.i_write | ~AESL_inst_myproject.layer7_out_60_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_60_V_U.i_write | ~AESL_inst_myproject.layer7_out_61_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_61_V_U.i_write | ~AESL_inst_myproject.layer7_out_62_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_62_V_U.i_write | ~AESL_inst_myproject.layer7_out_63_V_U.t_empty_n & (AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_ready | AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_63_V_U.i_write);
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_read);
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_read | ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_full_n & AESL_inst_myproject.clone_vec_ap_fixed_16_8_5_3_0_layer7_out_config_U0.ap_done & deadlock_detector.ap_done_reg_4 & ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[8 : 0] = dep_chan_data_4_5;
    assign token_in_vec_5[0] = token_4_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[17 : 9] = dep_chan_data_6_5;
    assign token_in_vec_5[1] = token_6_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_8_5;
    assign in_chan_dep_data_vec_5[26 : 18] = dep_chan_data_8_5;
    assign token_in_vec_5[2] = token_8_5;
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[0];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[1];
    assign dep_chan_vld_5_8 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_8 = out_chan_dep_data_5;
    assign token_5_8 = token_out_vec_5[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$edge_aggregate_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$edge_aggregate_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$edge_aggregate_U0$ap_idle <= AESL_inst_myproject.edge_aggregate_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.edge_aggregate_U0
    AESL_deadlock_detect_unit #(9, 6, 3, 3) AESL_deadlock_detect_unit_6 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (~AESL_inst_myproject.layer7_out_cpy1_0_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_0_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_1_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_2_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_3_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_4_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_5_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_6_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_7_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_8_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_9_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_10_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_11_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_12_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_13_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_14_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_15_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_16_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_17_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_18_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_19_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_20_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_21_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_22_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_23_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_24_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_25_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_26_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_27_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_28_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_29_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_30_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_31_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_32_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_33_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_34_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_35_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_36_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_37_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_38_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_39_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_40_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_41_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_42_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_43_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_44_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_45_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_46_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_47_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_48_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_49_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_50_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_51_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_52_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_53_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_54_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_55_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_56_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_57_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_58_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_59_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_60_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_61_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_62_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy1_63_V_U.i_write);
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (~AESL_inst_myproject.edge_index_cpy3_1_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_1_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_3_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_3_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_5_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_5_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_7_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_7_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_9_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_9_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_11_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_11_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_13_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_13_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_15_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_15_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_17_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_17_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_19_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_19_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_21_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_21_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_23_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_23_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_25_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_25_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_27_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_27_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_29_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_29_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy3_31_V_U.t_empty_n & (AESL_inst_myproject.edge_aggregate_U0.ap_ready | AESL_inst_myproject.edge_aggregate_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy3_31_V_U.i_write);
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (~AESL_inst_myproject.layer9_out_0_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_0_V_U.t_read | ~AESL_inst_myproject.layer9_out_1_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_1_V_U.t_read | ~AESL_inst_myproject.layer9_out_2_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_2_V_U.t_read | ~AESL_inst_myproject.layer9_out_3_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_3_V_U.t_read | ~AESL_inst_myproject.layer9_out_4_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_4_V_U.t_read | ~AESL_inst_myproject.layer9_out_5_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_5_V_U.t_read | ~AESL_inst_myproject.layer9_out_6_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_6_V_U.t_read | ~AESL_inst_myproject.layer9_out_7_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_7_V_U.t_read | ~AESL_inst_myproject.layer9_out_8_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_8_V_U.t_read | ~AESL_inst_myproject.layer9_out_9_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_9_V_U.t_read | ~AESL_inst_myproject.layer9_out_10_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_10_V_U.t_read | ~AESL_inst_myproject.layer9_out_11_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_11_V_U.t_read | ~AESL_inst_myproject.layer9_out_12_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_12_V_U.t_read | ~AESL_inst_myproject.layer9_out_13_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_13_V_U.t_read | ~AESL_inst_myproject.layer9_out_14_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_14_V_U.t_read | ~AESL_inst_myproject.layer9_out_15_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_15_V_U.t_read | ~AESL_inst_myproject.layer9_out_16_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_16_V_U.t_read | ~AESL_inst_myproject.layer9_out_17_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_17_V_U.t_read | ~AESL_inst_myproject.layer9_out_18_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_18_V_U.t_read | ~AESL_inst_myproject.layer9_out_19_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_19_V_U.t_read | ~AESL_inst_myproject.layer9_out_20_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_20_V_U.t_read | ~AESL_inst_myproject.layer9_out_21_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_21_V_U.t_read | ~AESL_inst_myproject.layer9_out_22_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_22_V_U.t_read | ~AESL_inst_myproject.layer9_out_23_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_23_V_U.t_read | ~AESL_inst_myproject.layer9_out_24_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_24_V_U.t_read | ~AESL_inst_myproject.layer9_out_25_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_25_V_U.t_read | ~AESL_inst_myproject.layer9_out_26_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_26_V_U.t_read | ~AESL_inst_myproject.layer9_out_27_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_27_V_U.t_read | ~AESL_inst_myproject.layer9_out_28_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_28_V_U.t_read | ~AESL_inst_myproject.layer9_out_29_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_29_V_U.t_read | ~AESL_inst_myproject.layer9_out_30_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_30_V_U.t_read | ~AESL_inst_myproject.layer9_out_31_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_31_V_U.t_read | ~AESL_inst_myproject.layer9_out_32_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_32_V_U.t_read | ~AESL_inst_myproject.layer9_out_33_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_33_V_U.t_read | ~AESL_inst_myproject.layer9_out_34_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_34_V_U.t_read | ~AESL_inst_myproject.layer9_out_35_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_35_V_U.t_read | ~AESL_inst_myproject.layer9_out_36_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_36_V_U.t_read | ~AESL_inst_myproject.layer9_out_37_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_37_V_U.t_read | ~AESL_inst_myproject.layer9_out_38_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_38_V_U.t_read | ~AESL_inst_myproject.layer9_out_39_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_39_V_U.t_read | ~AESL_inst_myproject.layer9_out_40_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_40_V_U.t_read | ~AESL_inst_myproject.layer9_out_41_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_41_V_U.t_read | ~AESL_inst_myproject.layer9_out_42_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_42_V_U.t_read | ~AESL_inst_myproject.layer9_out_43_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_43_V_U.t_read | ~AESL_inst_myproject.layer9_out_44_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_44_V_U.t_read | ~AESL_inst_myproject.layer9_out_45_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_45_V_U.t_read | ~AESL_inst_myproject.layer9_out_46_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_46_V_U.t_read | ~AESL_inst_myproject.layer9_out_47_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_47_V_U.t_read | ~AESL_inst_myproject.layer9_out_48_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_48_V_U.t_read | ~AESL_inst_myproject.layer9_out_49_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_49_V_U.t_read | ~AESL_inst_myproject.layer9_out_50_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_50_V_U.t_read | ~AESL_inst_myproject.layer9_out_51_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_51_V_U.t_read | ~AESL_inst_myproject.layer9_out_52_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_52_V_U.t_read | ~AESL_inst_myproject.layer9_out_53_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_53_V_U.t_read | ~AESL_inst_myproject.layer9_out_54_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_54_V_U.t_read | ~AESL_inst_myproject.layer9_out_55_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_55_V_U.t_read | ~AESL_inst_myproject.layer9_out_56_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_56_V_U.t_read | ~AESL_inst_myproject.layer9_out_57_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_57_V_U.t_read | ~AESL_inst_myproject.layer9_out_58_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_58_V_U.t_read | ~AESL_inst_myproject.layer9_out_59_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_59_V_U.t_read | ~AESL_inst_myproject.layer9_out_60_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_60_V_U.t_read | ~AESL_inst_myproject.layer9_out_61_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_61_V_U.t_read | ~AESL_inst_myproject.layer9_out_62_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_62_V_U.t_read | ~AESL_inst_myproject.layer9_out_63_V_U.i_full_n & AESL_inst_myproject.edge_aggregate_U0.ap_done & deadlock_detector.ap_done_reg_5 & ~AESL_inst_myproject.layer9_out_63_V_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_3_6;
    assign in_chan_dep_data_vec_6[8 : 0] = dep_chan_data_3_6;
    assign token_in_vec_6[0] = token_3_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[17 : 9] = dep_chan_data_5_6;
    assign token_in_vec_6[1] = token_5_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[26 : 18] = dep_chan_data_7_6;
    assign token_in_vec_6[2] = token_7_6;
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[0];
    assign dep_chan_vld_6_3 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_3 = out_chan_dep_data_6;
    assign token_6_3 = token_out_vec_6[1];
    assign dep_chan_vld_6_7 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_7 = out_chan_dep_data_6;
    assign token_6_7 = token_out_vec_6[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0$ap_idle <= AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0
    AESL_deadlock_detect_unit #(9, 7, 3, 3) AESL_deadlock_detect_unit_7 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (~AESL_inst_myproject.node_attr_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_0_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_1_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_2_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_3_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_4_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_5_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_6_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_7_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_8_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_9_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_10_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_11_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_12_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_13_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_14_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_15_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_16_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_17_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_18_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_19_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_20_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_21_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_22_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_23_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_24_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_25_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_26_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_27_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_28_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_29_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_30_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_31_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_32_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_32_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_33_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_33_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_34_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_34_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_35_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_35_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_36_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_36_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_37_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_37_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_38_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_38_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_39_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_39_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_40_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_40_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_41_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_41_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_42_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_42_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_43_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_43_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_44_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_44_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_45_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_45_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_46_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_46_V_U.i_write | ~AESL_inst_myproject.node_attr_cpy2_47_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.node_attr_cpy2_47_V_U.i_write);
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (~AESL_inst_myproject.layer9_out_0_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_0_V_U.i_write | ~AESL_inst_myproject.layer9_out_1_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_1_V_U.i_write | ~AESL_inst_myproject.layer9_out_2_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_2_V_U.i_write | ~AESL_inst_myproject.layer9_out_3_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_3_V_U.i_write | ~AESL_inst_myproject.layer9_out_4_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_4_V_U.i_write | ~AESL_inst_myproject.layer9_out_5_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_5_V_U.i_write | ~AESL_inst_myproject.layer9_out_6_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_6_V_U.i_write | ~AESL_inst_myproject.layer9_out_7_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_7_V_U.i_write | ~AESL_inst_myproject.layer9_out_8_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_8_V_U.i_write | ~AESL_inst_myproject.layer9_out_9_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_9_V_U.i_write | ~AESL_inst_myproject.layer9_out_10_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_10_V_U.i_write | ~AESL_inst_myproject.layer9_out_11_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_11_V_U.i_write | ~AESL_inst_myproject.layer9_out_12_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_12_V_U.i_write | ~AESL_inst_myproject.layer9_out_13_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_13_V_U.i_write | ~AESL_inst_myproject.layer9_out_14_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_14_V_U.i_write | ~AESL_inst_myproject.layer9_out_15_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_15_V_U.i_write | ~AESL_inst_myproject.layer9_out_16_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_16_V_U.i_write | ~AESL_inst_myproject.layer9_out_17_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_17_V_U.i_write | ~AESL_inst_myproject.layer9_out_18_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_18_V_U.i_write | ~AESL_inst_myproject.layer9_out_19_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_19_V_U.i_write | ~AESL_inst_myproject.layer9_out_20_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_20_V_U.i_write | ~AESL_inst_myproject.layer9_out_21_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_21_V_U.i_write | ~AESL_inst_myproject.layer9_out_22_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_22_V_U.i_write | ~AESL_inst_myproject.layer9_out_23_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_23_V_U.i_write | ~AESL_inst_myproject.layer9_out_24_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_24_V_U.i_write | ~AESL_inst_myproject.layer9_out_25_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_25_V_U.i_write | ~AESL_inst_myproject.layer9_out_26_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_26_V_U.i_write | ~AESL_inst_myproject.layer9_out_27_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_27_V_U.i_write | ~AESL_inst_myproject.layer9_out_28_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_28_V_U.i_write | ~AESL_inst_myproject.layer9_out_29_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_29_V_U.i_write | ~AESL_inst_myproject.layer9_out_30_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_30_V_U.i_write | ~AESL_inst_myproject.layer9_out_31_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_31_V_U.i_write | ~AESL_inst_myproject.layer9_out_32_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_32_V_U.i_write | ~AESL_inst_myproject.layer9_out_33_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_33_V_U.i_write | ~AESL_inst_myproject.layer9_out_34_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_34_V_U.i_write | ~AESL_inst_myproject.layer9_out_35_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_35_V_U.i_write | ~AESL_inst_myproject.layer9_out_36_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_36_V_U.i_write | ~AESL_inst_myproject.layer9_out_37_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_37_V_U.i_write | ~AESL_inst_myproject.layer9_out_38_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_38_V_U.i_write | ~AESL_inst_myproject.layer9_out_39_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_39_V_U.i_write | ~AESL_inst_myproject.layer9_out_40_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_40_V_U.i_write | ~AESL_inst_myproject.layer9_out_41_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_41_V_U.i_write | ~AESL_inst_myproject.layer9_out_42_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_42_V_U.i_write | ~AESL_inst_myproject.layer9_out_43_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_43_V_U.i_write | ~AESL_inst_myproject.layer9_out_44_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_44_V_U.i_write | ~AESL_inst_myproject.layer9_out_45_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_45_V_U.i_write | ~AESL_inst_myproject.layer9_out_46_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_46_V_U.i_write | ~AESL_inst_myproject.layer9_out_47_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_47_V_U.i_write | ~AESL_inst_myproject.layer9_out_48_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_48_V_U.i_write | ~AESL_inst_myproject.layer9_out_49_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_49_V_U.i_write | ~AESL_inst_myproject.layer9_out_50_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_50_V_U.i_write | ~AESL_inst_myproject.layer9_out_51_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_51_V_U.i_write | ~AESL_inst_myproject.layer9_out_52_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_52_V_U.i_write | ~AESL_inst_myproject.layer9_out_53_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_53_V_U.i_write | ~AESL_inst_myproject.layer9_out_54_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_54_V_U.i_write | ~AESL_inst_myproject.layer9_out_55_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_55_V_U.i_write | ~AESL_inst_myproject.layer9_out_56_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_56_V_U.i_write | ~AESL_inst_myproject.layer9_out_57_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_57_V_U.i_write | ~AESL_inst_myproject.layer9_out_58_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_58_V_U.i_write | ~AESL_inst_myproject.layer9_out_59_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_59_V_U.i_write | ~AESL_inst_myproject.layer9_out_60_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_60_V_U.i_write | ~AESL_inst_myproject.layer9_out_61_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_61_V_U.i_write | ~AESL_inst_myproject.layer9_out_62_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_62_V_U.i_write | ~AESL_inst_myproject.layer9_out_63_V_U.t_empty_n & (AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_ready | AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_idle) & ~AESL_inst_myproject.layer9_out_63_V_U.i_write);
    assign proc_dep_vld_vec_7[2] = dl_detect_out ? proc_dep_vld_vec_7_reg[2] : (~AESL_inst_myproject.layer10_out_0_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_0_V_U.t_read | ~AESL_inst_myproject.layer10_out_1_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_1_V_U.t_read | ~AESL_inst_myproject.layer10_out_2_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_2_V_U.t_read | ~AESL_inst_myproject.layer10_out_3_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_3_V_U.t_read | ~AESL_inst_myproject.layer10_out_4_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_4_V_U.t_read | ~AESL_inst_myproject.layer10_out_5_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_5_V_U.t_read | ~AESL_inst_myproject.layer10_out_6_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_6_V_U.t_read | ~AESL_inst_myproject.layer10_out_7_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_7_V_U.t_read | ~AESL_inst_myproject.layer10_out_8_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_8_V_U.t_read | ~AESL_inst_myproject.layer10_out_9_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_9_V_U.t_read | ~AESL_inst_myproject.layer10_out_10_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_10_V_U.t_read | ~AESL_inst_myproject.layer10_out_11_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_11_V_U.t_read | ~AESL_inst_myproject.layer10_out_12_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_12_V_U.t_read | ~AESL_inst_myproject.layer10_out_13_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_13_V_U.t_read | ~AESL_inst_myproject.layer10_out_14_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_14_V_U.t_read | ~AESL_inst_myproject.layer10_out_15_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_15_V_U.t_read | ~AESL_inst_myproject.layer10_out_16_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_16_V_U.t_read | ~AESL_inst_myproject.layer10_out_17_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_17_V_U.t_read | ~AESL_inst_myproject.layer10_out_18_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_18_V_U.t_read | ~AESL_inst_myproject.layer10_out_19_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_19_V_U.t_read | ~AESL_inst_myproject.layer10_out_20_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_20_V_U.t_read | ~AESL_inst_myproject.layer10_out_21_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_21_V_U.t_read | ~AESL_inst_myproject.layer10_out_22_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_22_V_U.t_read | ~AESL_inst_myproject.layer10_out_23_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_23_V_U.t_read | ~AESL_inst_myproject.layer10_out_24_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_24_V_U.t_read | ~AESL_inst_myproject.layer10_out_25_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_25_V_U.t_read | ~AESL_inst_myproject.layer10_out_26_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_26_V_U.t_read | ~AESL_inst_myproject.layer10_out_27_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_27_V_U.t_read | ~AESL_inst_myproject.layer10_out_28_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_28_V_U.t_read | ~AESL_inst_myproject.layer10_out_29_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_29_V_U.t_read | ~AESL_inst_myproject.layer10_out_30_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_30_V_U.t_read | ~AESL_inst_myproject.layer10_out_31_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_31_V_U.t_read | ~AESL_inst_myproject.layer10_out_32_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_32_V_U.t_read | ~AESL_inst_myproject.layer10_out_33_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_33_V_U.t_read | ~AESL_inst_myproject.layer10_out_34_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_34_V_U.t_read | ~AESL_inst_myproject.layer10_out_35_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_35_V_U.t_read | ~AESL_inst_myproject.layer10_out_36_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_36_V_U.t_read | ~AESL_inst_myproject.layer10_out_37_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_37_V_U.t_read | ~AESL_inst_myproject.layer10_out_38_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_38_V_U.t_read | ~AESL_inst_myproject.layer10_out_39_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_39_V_U.t_read | ~AESL_inst_myproject.layer10_out_40_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_40_V_U.t_read | ~AESL_inst_myproject.layer10_out_41_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_41_V_U.t_read | ~AESL_inst_myproject.layer10_out_42_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_42_V_U.t_read | ~AESL_inst_myproject.layer10_out_43_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_43_V_U.t_read | ~AESL_inst_myproject.layer10_out_44_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_44_V_U.t_read | ~AESL_inst_myproject.layer10_out_45_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_45_V_U.t_read | ~AESL_inst_myproject.layer10_out_46_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_46_V_U.t_read | ~AESL_inst_myproject.layer10_out_47_V_U.i_full_n & AESL_inst_myproject.nodeblock_ap_fixed_ap_fixed_16_8_5_3_0_config10_U0.ap_done & deadlock_detector.ap_done_reg_6 & ~AESL_inst_myproject.layer10_out_47_V_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_1_7;
    assign in_chan_dep_data_vec_7[8 : 0] = dep_chan_data_1_7;
    assign token_in_vec_7[0] = token_1_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_6_7;
    assign in_chan_dep_data_vec_7[17 : 9] = dep_chan_data_6_7;
    assign token_in_vec_7[1] = token_6_7;
    assign in_chan_dep_vld_vec_7[2] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[26 : 18] = dep_chan_data_8_7;
    assign token_in_vec_7[2] = token_8_7;
    assign dep_chan_vld_7_1 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_1 = out_chan_dep_data_7;
    assign token_7_1 = token_out_vec_7[0];
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[1];
    assign dep_chan_vld_7_8 = out_chan_dep_vld_vec_7[2];
    assign dep_chan_data_7_8 = out_chan_dep_data_7;
    assign token_7_8 = token_out_vec_7[2];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myproject$edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0$ap_idle <= AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0
    AESL_deadlock_detect_unit #(9, 8, 3, 3) AESL_deadlock_detect_unit_8 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (~AESL_inst_myproject.layer10_out_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_0_V_U.i_write | ~AESL_inst_myproject.layer10_out_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_1_V_U.i_write | ~AESL_inst_myproject.layer10_out_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_2_V_U.i_write | ~AESL_inst_myproject.layer10_out_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_3_V_U.i_write | ~AESL_inst_myproject.layer10_out_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_4_V_U.i_write | ~AESL_inst_myproject.layer10_out_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_5_V_U.i_write | ~AESL_inst_myproject.layer10_out_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_6_V_U.i_write | ~AESL_inst_myproject.layer10_out_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_7_V_U.i_write | ~AESL_inst_myproject.layer10_out_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_8_V_U.i_write | ~AESL_inst_myproject.layer10_out_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_9_V_U.i_write | ~AESL_inst_myproject.layer10_out_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_10_V_U.i_write | ~AESL_inst_myproject.layer10_out_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_11_V_U.i_write | ~AESL_inst_myproject.layer10_out_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_12_V_U.i_write | ~AESL_inst_myproject.layer10_out_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_13_V_U.i_write | ~AESL_inst_myproject.layer10_out_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_14_V_U.i_write | ~AESL_inst_myproject.layer10_out_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_15_V_U.i_write | ~AESL_inst_myproject.layer10_out_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_16_V_U.i_write | ~AESL_inst_myproject.layer10_out_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_17_V_U.i_write | ~AESL_inst_myproject.layer10_out_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_18_V_U.i_write | ~AESL_inst_myproject.layer10_out_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_19_V_U.i_write | ~AESL_inst_myproject.layer10_out_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_20_V_U.i_write | ~AESL_inst_myproject.layer10_out_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_21_V_U.i_write | ~AESL_inst_myproject.layer10_out_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_22_V_U.i_write | ~AESL_inst_myproject.layer10_out_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_23_V_U.i_write | ~AESL_inst_myproject.layer10_out_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_24_V_U.i_write | ~AESL_inst_myproject.layer10_out_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_25_V_U.i_write | ~AESL_inst_myproject.layer10_out_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_26_V_U.i_write | ~AESL_inst_myproject.layer10_out_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_27_V_U.i_write | ~AESL_inst_myproject.layer10_out_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_28_V_U.i_write | ~AESL_inst_myproject.layer10_out_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_29_V_U.i_write | ~AESL_inst_myproject.layer10_out_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_30_V_U.i_write | ~AESL_inst_myproject.layer10_out_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_31_V_U.i_write | ~AESL_inst_myproject.layer10_out_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_32_V_U.i_write | ~AESL_inst_myproject.layer10_out_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_33_V_U.i_write | ~AESL_inst_myproject.layer10_out_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_34_V_U.i_write | ~AESL_inst_myproject.layer10_out_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_35_V_U.i_write | ~AESL_inst_myproject.layer10_out_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_36_V_U.i_write | ~AESL_inst_myproject.layer10_out_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_37_V_U.i_write | ~AESL_inst_myproject.layer10_out_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_38_V_U.i_write | ~AESL_inst_myproject.layer10_out_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_39_V_U.i_write | ~AESL_inst_myproject.layer10_out_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_40_V_U.i_write | ~AESL_inst_myproject.layer10_out_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_41_V_U.i_write | ~AESL_inst_myproject.layer10_out_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_42_V_U.i_write | ~AESL_inst_myproject.layer10_out_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_43_V_U.i_write | ~AESL_inst_myproject.layer10_out_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_44_V_U.i_write | ~AESL_inst_myproject.layer10_out_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_45_V_U.i_write | ~AESL_inst_myproject.layer10_out_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_46_V_U.i_write | ~AESL_inst_myproject.layer10_out_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer10_out_47_V_U.i_write);
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (~AESL_inst_myproject.layer7_out_cpy2_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_0_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_1_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_2_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_3_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_4_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_5_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_6_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_7_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_8_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_9_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_10_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_11_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_12_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_13_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_14_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_15_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_16_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_17_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_18_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_19_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_20_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_21_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_22_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_23_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_24_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_25_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_26_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_27_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_28_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_29_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_30_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_31_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_32_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_33_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_34_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_35_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_36_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_37_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_38_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_39_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_40_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_41_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_42_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_43_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_44_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_45_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_46_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_47_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_48_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_49_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_50_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_51_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_52_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_53_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_54_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_55_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_56_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_57_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_58_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_59_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_60_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_61_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_62_V_U.i_write | ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.layer7_out_cpy2_63_V_U.i_write);
    assign proc_dep_vld_vec_8[2] = dl_detect_out ? proc_dep_vld_vec_8_reg[2] : (~AESL_inst_myproject.edge_index_cpy4_0_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_0_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_1_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_1_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_2_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_2_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_3_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_3_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_4_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_4_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_5_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_5_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_6_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_6_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_7_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_7_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_8_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_8_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_9_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_9_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_10_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_10_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_11_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_11_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_12_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_12_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_13_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_13_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_14_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_14_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_15_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_15_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_16_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_16_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_17_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_17_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_18_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_18_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_19_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_19_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_20_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_20_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_21_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_21_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_22_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_22_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_23_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_23_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_24_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_24_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_25_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_25_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_26_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_26_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_27_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_27_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_28_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_28_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_29_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_29_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_30_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_30_V_U.i_write | ~AESL_inst_myproject.edge_index_cpy4_31_V_U.t_empty_n & (AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_ready | AESL_inst_myproject.edgeblock_ap_fixed_ap_uint_ap_fixed_config11_U0.ap_idle) & ~AESL_inst_myproject.edge_index_cpy4_31_V_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_3_8;
    assign in_chan_dep_data_vec_8[8 : 0] = dep_chan_data_3_8;
    assign token_in_vec_8[0] = token_3_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_5_8;
    assign in_chan_dep_data_vec_8[17 : 9] = dep_chan_data_5_8;
    assign token_in_vec_8[1] = token_5_8;
    assign in_chan_dep_vld_vec_8[2] = dep_chan_vld_7_8;
    assign in_chan_dep_data_vec_8[26 : 18] = dep_chan_data_7_8;
    assign token_in_vec_8[2] = token_7_8;
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[0];
    assign dep_chan_vld_8_5 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_5 = out_chan_dep_data_8;
    assign token_8_5 = token_out_vec_8[1];
    assign dep_chan_vld_8_3 = out_chan_dep_vld_vec_8[2];
    assign dep_chan_data_8_3 = out_chan_dep_data_8;
    assign token_8_3 = token_out_vec_8[2];


    AESL_deadlock_report_unit #(9) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
